package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "../AXI_Lite_UVM_Agent/src/axi_lite_include.svh"
    `include "axi_lite_cnt_sequence_config.svh"
    `include "axi_lite_cnt_sequence.svh"
    `include "test_env.svh"
    `include "base_test.svh"
    
endpackage